library verilog;
use verilog.vl_types.all;
entity arith_tb is
end arith_tb;
