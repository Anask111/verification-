library verilog;
use verilog.vl_types.all;
entity fact_test is
end fact_test;
