library verilog;
use verilog.vl_types.all;
entity fifo_tb1 is
end fifo_tb1;
