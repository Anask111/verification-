library verilog;
use verilog.vl_types.all;
entity and1_tb is
end and1_tb;
