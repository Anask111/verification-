library verilog;
use verilog.vl_types.all;
entity HAcase_tb is
end HAcase_tb;
