library verilog;
use verilog.vl_types.all;
entity que is
end que;
