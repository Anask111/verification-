library verilog;
use verilog.vl_types.all;
entity nand1_tb is
end nand1_tb;
