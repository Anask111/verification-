library verilog;
use verilog.vl_types.all;
entity decoderc_tb is
end decoderc_tb;
