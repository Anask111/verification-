library verilog;
use verilog.vl_types.all;
entity odd_tb is
end odd_tb;
