//module muxr4 (y,a,b,c,d,s1,s2,s3);
//output  y;
//input [7:0] a,b,c,d;
//input [4:0]s;
//
//
////assign y = s1?(s0:d:c):(s0?b:a);
//// 8:1 mux
// (s[4]?
//   (s[3]?( 
//	   s[2]?( s[1]?(((s[0]?a[0]:a[1]):(s[0]?a[2]:a[3])):(s[0]?a[4]:a[5]):(s[0]?a[6]:a[7]))):((s[0]?b[0]:b[1]):(s[0]?b[2]:b[3])):(s[0]?b[4]:b[5]):(s[0]?b[6]:b[7]))))):( s[1]?(((s[0]?c[0]:c[1]):(s[0]?c[2]:c[3])):(s[0]?(c[4]:c[5]):(s[0]?c[6]:c[7]))) :((s[0]?d[0]:d[1]):(s[0]?d[2]:d[3])):(s[0]?(d[4]:d[5]):(s[0]?d[6]:d[7])))))) 
//		:( s[2]?( s[1]?(((s[0]?a[0]:a[1]):(s[0]?a[2]:a[3])):(s[0]?a[4]:a[5]):(s[0]?a[6]:a[7]))) :((s[0]?b[0]:b[1]):(s[0]?b[2]:b[3])):(s[0]?(b[4]:b[5]):(s[0]?b[6]:b[7]))))) :( s[1]?(((s[0]?c[0]:c[1]):(s[0]?c[2]:c[3])):(s[0]?c[4]:c[5]):(s[0]?c[6]:c[7]))) :((s[0]?d[0]:d[1]):(s[0]?d[2]:d[3])):(s[0]?d[4]:d[5]):(s[0]?d[6]:d[7])))))))
//	 :(s[3]?( s[2]?( s[1]?(((s[0]?a[0]:a[1]):(s[0]?a[2]:a[3])):(s[0]?a[4]:a[5]):(s[0]?a[6]:a[7]))) :((s[0]?b[0]:b[1]):(s[0]?b[2]:b[3])):(s[0]?b[4]:b[5]):(s[0]?b[6]:b[7]))))):( s[1]?(((s[0]?c[0]:c[1]):(s[0]?c[2]:c[3])):(s[0]?c[4]:c[5]):(s[0]?c[6]:c[7]))) :((s[0]?d[0]:d[1]):(s[0]?d[2]:d[3])):(s[0]?(d[4]:d[5]):(s[0]?d[6]:d[7])))))) 
//	   :( s[2]?( s[1]?(((s[0]?a[0]:a[1]):(s[0]?a[2]:a[3])):(s[0]?(a[4]:a[5]):(s[0]?a[6]:a[7]))) :((s[0]?b[0]:b[1]):(s[0]?b[2]:b[3])):(s[0]?b[4]:b[5]):(s[0]?b[6]:b[7]))))) :( s[1]?(((s[0]?c[0]:c[1]):(s[0]?c[2]:c[3])):(s[0]?c[4]:c[5]):(s[0]?c[6]:c[7]))) :((s[0]?d[0]:d[1]):(s[0]?d[2]:d[3])):(s[0]?d[4]:d[5]):(s[0]?d[6]:d[7]))))))))	
//			 
//endmodule


module muxr4_tb;
  reg s1,s2;
  reg a,b,c,d;
  wire y;
  muxr4 i_muxr4(y,a,b,c,d,s1,s2);
 
  initial
  begin
  $monitor("At time %0t - a=%b, b=%b ,c=%b, d=%b , y=%b,s1=%b,s2=%b ",$time,y,a,b,c,d,s1,s2);
  a ='b1;
  b='b1;
  c ='b1;
  d='b1;
  s1='b1;
  s2='b0;
end

   always #1 a=~a;
  always #2 b=~b;
 always #3 c=~c;
  always #4 d=~d;
   always #5 s1=~s1;
always #10 s2=~s2;

initial #200$finish;
endmodule
