library verilog;
use verilog.vl_types.all;
entity sumdif_tb is
end sumdif_tb;
