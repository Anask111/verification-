library verilog;
use verilog.vl_types.all;
entity hadder_tb is
end hadder_tb;
