library verilog;
use verilog.vl_types.all;
entity dl_tb is
end dl_tb;
