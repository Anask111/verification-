library verilog;
use verilog.vl_types.all;
entity bintogre_tb is
end bintogre_tb;
