library verilog;
use verilog.vl_types.all;
entity ANDtb is
end ANDtb;
