library verilog;
use verilog.vl_types.all;
entity reverse_test is
end reverse_test;
