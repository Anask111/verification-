library verilog;
use verilog.vl_types.all;
entity muxr_tb is
end muxr_tb;
