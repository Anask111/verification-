library verilog;
use verilog.vl_types.all;
entity compr2_tb is
end compr2_tb;
