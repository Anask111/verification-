library verilog;
use verilog.vl_types.all;
entity mealy1010na_tb is
end mealy1010na_tb;
