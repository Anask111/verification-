library verilog;
use verilog.vl_types.all;
entity greytobin_tb is
end greytobin_tb;
