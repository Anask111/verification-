library verilog;
use verilog.vl_types.all;
entity demux_tb is
end demux_tb;
