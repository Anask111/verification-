library verilog;
use verilog.vl_types.all;
entity FA_tb is
end FA_tb;
