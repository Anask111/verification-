library verilog;
use verilog.vl_types.all;
entity mealy1010a_tb is
end mealy1010a_tb;
