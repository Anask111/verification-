library verilog;
use verilog.vl_types.all;
entity moore1010na_tb is
end moore1010na_tb;
