library verilog;
use verilog.vl_types.all;
entity demuxc_tb is
end demuxc_tb;
