library verilog;
use verilog.vl_types.all;
entity moore1010a_tb is
end moore1010a_tb;
