library verilog;
use verilog.vl_types.all;
entity file_write is
end file_write;
