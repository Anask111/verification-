library verilog;
use verilog.vl_types.all;
entity comp2_tb is
end comp2_tb;
