library verilog;
use verilog.vl_types.all;
entity xnor1_tb is
end xnor1_tb;
