library verilog;
use verilog.vl_types.all;
entity seven_TB is
end seven_TB;
