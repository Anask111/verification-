library verilog;
use verilog.vl_types.all;
entity duty_tb is
end duty_tb;
