library verilog;
use verilog.vl_types.all;
entity sr_tb is
end sr_tb;
