library verilog;
use verilog.vl_types.all;
entity ORtb is
end ORtb;
