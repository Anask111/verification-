library verilog;
use verilog.vl_types.all;
entity nor1_tb is
end nor1_tb;
