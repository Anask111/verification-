library verilog;
use verilog.vl_types.all;
entity HA_tb is
end HA_tb;
