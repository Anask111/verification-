library verilog;
use verilog.vl_types.all;
entity inv is
    port(
        \out\           : out    vl_logic;
        \in\            : in     vl_logic
    );
end inv;
