library verilog;
use verilog.vl_types.all;
entity rough_sv_unit is
end rough_sv_unit;
