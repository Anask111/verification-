library verilog;
use verilog.vl_types.all;
entity arrtb is
end arrtb;
