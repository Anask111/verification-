library verilog;
use verilog.vl_types.all;
entity xor1_tb is
end xor1_tb;
