library verilog;
use verilog.vl_types.all;
entity fa_tb is
end fa_tb;
