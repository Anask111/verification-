library verilog;
use verilog.vl_types.all;
entity file_read is
end file_read;
