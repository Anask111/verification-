library verilog;
use verilog.vl_types.all;
entity oddp_tb is
end oddp_tb;
