library verilog;
use verilog.vl_types.all;
entity xnor1 is
    port(
        \out\           : out    vl_logic;
        in1             : in     vl_logic;
        in2             : in     vl_logic
    );
end xnor1;
