library verilog;
use verilog.vl_types.all;
entity bintogrey_tb is
end bintogrey_tb;
