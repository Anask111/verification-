library verilog;
use verilog.vl_types.all;
entity JK_tb is
end JK_tb;
