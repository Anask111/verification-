library verilog;
use verilog.vl_types.all;
entity encoder8_tb is
end encoder8_tb;
