library verilog;
use verilog.vl_types.all;
entity muxr4_tb is
end muxr4_tb;
