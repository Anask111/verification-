library verilog;
use verilog.vl_types.all;
entity or1_tb is
end or1_tb;
