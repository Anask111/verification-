library verilog;
use verilog.vl_types.all;
entity FAcase_tb is
end FAcase_tb;
