library verilog;
use verilog.vl_types.all;
entity fig1_tb is
end fig1_tb;
